SV_WU#0
SV_LF#0
SV_CR#0
SV_CG#0
SV_CL#0
SV_AK#0
LS_CR#0
LS_CL#0
LS_CG#0